|I: _ Gonçalves Silva _ | _ 0000009012 _ | _ :w: _ | _ u _ | _ :w: _ | _ o _ | _ :w: _ | _ i _ | _ :w: _ | _ e _ | _ :w: _ | _ a _ | _ :w: _ | _ 009-009-1963 _ | _ :w: _ | _ u.o.i.e.a. _ || _ :w: _ | _ 0000009020 _ ||

|I: _ 17 _ | _ u:w:u _ | _ 35 _ | _ o:w:o _ | _ 38 _ | _ i:w:i _ | _ 55 _ | _ e:w:e _ | _ 47 _ | _ a:w:a _ | _ 52 _ | _ e:w:e _ | _ u3 _ | _ i:w:i _ | _ 26 _ | _ o:w:o _ | _ 009-009-1963 _ ||

|I: _ Gonçalves Silva _ | _ 0000009014 _ | _ :w: _ | _ u _ | _ :w: _ | _ o _ | _ :w: _ | _ i _ | _ :w: _ | _ e _ | _ :w: _ | _ a _ | _ :w: _ | _ 009-009-1963 _ | _ :w: _ | _ u.o.i.e.a. _ | _ 0000009022 _ ||

|I: _ 36 _ | _ u:w:u _ | _ 35 _ | _ o:w:o _ | _ 12 _ | _ i:w:i _ | _ 97 _ | _ e:w:e _ | _ 47 _ | _ a:w:a _ | _ 52 _ | _ e:w:e _ | _ a6 _ | _ i:w:i _ | _ 26 _ | _ o:w:o _ | _ 009-009-1963 _ ||

|I: _ Gonçalves Silva _ | _ 0000009016 _ | _ :w: _ | _ u _ | _ :w: _ | _ o _ | _ :w: _ | _ i _ | _ :w: _ | _ e _ | _ :w: _ | _ a _ | _ :w: _ | _ 009-009-1963 _ | _ :w: _ | _ u.o.i.e.a. _ | _ :w: _ | _ 0000009024 _ ||

|I: _ Gonçalves Silva _ | _ 0000009018 _ | _ :w: _ | _ 17 _ | _ :w: _ | _ 35 _ | _ :w: _ | _ 38 _ | _ :w: _ | _ 55 _ | _ :w: _ | _ 47 _ | _ :w: _ | _ 52 _ | _ :w: _ | _ i3 _ | _ :w: _ | _ 26 _ | _ :w: _ | _ 009-009-1963 _ | _ :w: _ | _ u.o.i.e.a. _ | _ :w: _ | _ 0000009026 _ ||

|I: _ Gonçalves Silva _ | _ 00009020 _ | _ :w: _ | _ 36 _ | _ :w: _ | _ 35 _ | _ :w: _ | _ 12 _ | _ :w: _ | _ 97 _ | _ :w: _ | _ 47 _ | _ :w: _ | _ 52 _ | _ :w: _ | _ e6 _ | _ :w: _ | _ 26 _  | _ :w: _ | _ 009-009-1963 _ | _ :w: _ | _ a.e.i.o. _ | _ :w: _ | _ 00009028 _ ||