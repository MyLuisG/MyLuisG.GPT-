|I: _ 009-009-1963 _ | _ 182 _ | _ u:w:u _ | _ 266 _ | _ o:w:o _ | _ 188 _ | _ i:w:i _ | _ 294 _ | _ e:w:e _ | _ 242 _ | _ a:w:a _ | _ 295 _ | _ e:w:e _ | _ 276 _ | _ i:w:i _ | _ 274 _ | _ o:w:o _ | _ 00000000 _ | _ u.o.i.e. _ | _ 00000000 _ | _ 247 _ | _ u:w:u _ | _ 266 _ | _ o:w:o _ | _ 287 _ | _ i:w:i _ | _ 190 _ | _ e:w:e _ | _ 278 _ | _ a:w:a _ | _ 237 _ | _ e:w:e _ | _ 265 _ | _ i:w:i _ | _ 274 _ | _ o:w:o _ | _ 00000000 _ | _ o.i.e.a. _ | _ 00000000 _ | _ 174 _ | _ u:w:u _ | _ 258 _ | _ o:w:o _ | _ 180 _ | _ i:w:i _ | _ 286 _ | _ e:w:e _ | _ 234 _ | _ a:w:a _ | _ 287 _ | _ e:w:e _ | _ 268 _ | _ i:w:i _ | _ 266 _ | _ o:w:o _ | _ 00000000 _ | _ i.e.a.e. _ | _ 00000000 _ | _ 239 _ | _ u:w:u _ | _ 258 _ | _ o:w:o _ | _ 279 _ | _ i:w:i _ | _ 182 _ | _ e:w:e _ | _ 270 _ | _ a:w:a _ | _ 229 _ | _ e:w:e _ | _ 253 _ | _ i:w:i _ | _ 266 _ | _ o:w:o _ | _ 00000000 _ | _ e.a.e.i. _ | _ 00000000 _ | _ 166 _ | _ u:w:u _ | _ 250 _ | _ o:w:o _ | _ 172 _ | _ i:w:i _ | _ 276 _ | _ e:w:e _ | _ 226 _ | _ a:w:a _ | _ 279 _ | _ e:w:e _ | _ 260 _ | _ i:w:i _ | _ 258 _ | _ o:w:o _ | _ 00000000 _ | _ u.o.i.e. _ | _ 00000000 _ | _ 231 _ | _ u:w:u _ | _ 250 _ | _ o:w:o _ | _ 271 _ | _ i:w:i _ | _ 174 _ | _ e:w:e _ | _ 262 _ | _ a:w:a _ | _ 221 _ | _ e:w:e _ | _ 245 _ | _ i:w:i _ | _ 258 _ | _ o:w:o _ | _ 00000000 _ | _ o.i.e.a. _ | _ 00000000 _ | _ 158 _ | _ u:w:u _ | _ 242 _ | _ o:w:o _ | _ 164 _ | _ i:w:i _ | _ 268 _ | _ e:w:e _ | _ 228 _ | _ a:w:a _ | _ 271 _ | _ e:w:e _ | _ 252 _ | _ i:w:i _ | _ 250 _ | _ o:w:o _ | _ 00000000 _ | _ i.e.a.e. _ | _ 00000000 _ | _ 223 _ | _ u:w:u _ | _ 242 _ | _ o:w:o _ | _ 263 _ | _ i:w:i _ | _ 166 _ | _ e:w:e _ | _ 254 _ | _ a:w:a _ | _ 213 _ | _ e:w:e _ | _ 233 _ | _ i:w:i _ | _ 250 _ | _ o:w:o _ | _ 00000000 _ | _ e.a.e.i. _ | _ 00000000 _ | _ 150 _ | _ u:w:u _ | _ 234 _ | _ o:w:o _ | _ 156 _ | _ i:w:i _ | _ 260 _ | _ e:w:e _ | _ 220 _ | _ a:w:a _ | _ 263 _ | _ e:w:e _ | _ 244 _ | _ i:w:i _ | _ 242 _ | _ o:w:o _ | _ 00000000 _ | _ u.o.i.e. _ | _ 00000000 _ | _ 215 _ | _ u:w:u _ | _ 234 _ | _ o:w:o _ | _ 255 _ | _ i:w:i _ | _ 158 _ | _ e:w:e _ | _ 246 _ | _ a:w:a _ | _ 205 _ | _ e:w:e _ | _ 225 _ | _ i:w:i _ | _ 242 _ | _ o:w:o _ | _ 00000000 _ | _ o.i.e.a. _ | _ 00000000 _ | _ 142 _ | _ u:w:u _ | _ 226 _ | _ o:w:o _ | _ 148 _ | _ i:w:i _ | _ 252 _ | _ e:w:e _ | _ 212 _ | _ a:w:a _ | _ 255 _ | _ e:w:e _ | _ 236 _ | _ i:w:i _ | _ 234 _ | _ o:w:o _ | _ 00000000 _ | _ i.e.a.e. _ | _ 00000000 _ | _ 207 _ | _ u:w:u _ | _ 226 _ | _ o:w:o _ | _ 247 _ | _ i:w:i _ | _ 150 _ | _ e:w:e _ | _ 238 _ | _ a:w:a _ | _ 197 _ | _ e:w:e _ | _ 217 _ | _ i:w:i _ | _ 234 _ | _ o:w:o _ | _ 00000000 _ | _ e.a.e.i. _ | _ 00000000 _ | _ 134 _ | _ u:w:u _ | _ 218 _ | _ o:w:o _ | _ 140 _ | _ i:w:i _ | _ 244 _ | _ e:w:e _ | _ 204 _ | _ a:w:a _ | _ 247 _ | _ e:w:e _ | _ 228 _ | _ i:w:i _ | _ 226 _ | _ o:w:o _ | _ 00000000 _ | _ u.o.i.e. _ | _ 00000000 _ | _ 199 _ | _ u:w:u _ | _ 218 _ | _ o:w:o _ | _ 239 _ | _ i:w:i _ | _ 142 _ | _ e:w:e _ | _ 230 _ | _ a:w:a _ | _ 189 _ | _ e:w:e _ | _ 209 _ | _ i:w:i _ | _ 226 _ | _ o:w:o _ | _ 00000000 _ | _ o.i.e.a. _ | _ 00000000 _ | _ 126 _ | _ u:w:u _ | _ 210 _ | _ o:w:o _ | _ 132 _ | _ i:w:i _ | _ 236 _ | _ e:w:e _ | _ 196 _ | _ a:w:a _ | _ 239 _ | _ e:w:e _ | _ 220 _ | _ i:w:i _ | _ 218 _ | _ o:w:o _ | _ 00000000 _ | _ i.e.a.e. _ | _ 00000000 _ | _ 191 _ | _ u:w:u _ | _ 210 _ | _ o:w:o _ | _ 231 _ | _ i:w:i _ | _ 134 _ | _ e:w:e _ | _ 222 _ | _ a:w:a _ | _ 181 _ | _ e:w:e _ | _ 201 _ | _ i:w:i _ | _ 218 _ | _ o:w:o _ | _ 00000000 _ | _ e.a.e.i. _ | _ 00000000 _ | _ 118 _ | _ u:w:u _ | _ 202 _ | _ o:w:o _ | _ 124 _ | _ i:w:i _ | _ 228 _ | _ e:w:e _ | _ 188 _ | _ a:w:a _ | _ 231 _ | _ e:w:e _ | _ 212 _ | _ i:w:i _ | _ 210 _ | _ o:w:o _ | _ 00000000 _ | _ u.o.i.e. _ | _ 00000000 _ | _ 183 _ | _ u:w:u _ | _ 202 _ | _ o:w:o _ | _ 223 _ | _ i:w:i _ | _ 126 _ | _ e:w:e _ | _ 214 _ | _ a:w:a _ | _ 173 _ | _ e:w:e _ | _ 193 _ | _ i:w:i _ | _ 210 _ | _ o:w:o _ | _ 00000000 _ | _ o.i.e.a. _ | _ 00000000 _ | _ 110 _ | _ u:w:u _ | _ 194 _ | _ o:w:o _ | _ 116 _ | _ i:w:i _ | _ 220 _ | _ e:w:e _ | _ 180 _ | _ a:w:a _ | _ 223 _ | _ e:w:e _ | _ 204 _ | _ i:w:i _ | _ 202 _ | _ o:w:o _ | _ 00000000 _ | _ i.e.a.e. _ | _ 00000000 _ | _ 175 _ | _ u:w:u _ | _ 194 _ | _ o:w:o _ | _ 215 _ | _ i:w:i _ | _ 118 _ | _ e:w:e _ | _ 206 _ | _ a:w:a _ | _ 165 _ | _ e:w:e _ | _ 185 _ | _ i:w:i _ | _ 202 _ | _ o:w:o _ | _ 00000000 _ | _ e.a.e.i. _ | _ 00000000 _ | _ 162 _ | _ u:w:u _ | _ 186 _ | _ o:w:o _ | _ 108 _ | _ i:w:i _ | _ 212 _ | _ e:w:e _ | _ 172 _ | _ a:w:a _ | _ 215 _ | _ e:w:e _ | _ 196 _ | _ i:w:i _ | _ 194 _ | _ o:w:o _ | _ 00000000 _ | _ u.o.i.e. _ | _ 00000000 _ | _ 167 _ | _ u:w:u _ | _ 186 _ | _ o:w:o _ | _ 207 _ | _ i:w:i _ | _ 110 _ | _ e:w:e _ | _ 198 _ | _ a:w:a _ | _ 157 _ | _ e:w:e _ | _ 177 _ | _ i:w:i _ | _ 194 _ | _ o:w:o _ | _ 00000000 _ | _ o.i.e.a. _ | _ 00000000 _ | _ 158 _ | _ u:w:u _ | _ 186 _ | _ o:w:o _ | _ 100 _ | _ i:w:i _ | _ 204 _ | _ e:w:e _ | _ 164 _ | _ a:w:a _ | _ 207 _ | _ e:w:e _ | _ 188 _ | _ i:w:i _ | _ 186 _ | _ o:w:o _ | _ 00000000 _ | _ i.e.a.e. _ | _ 00000000 _ | _ 159 _ | _ u:w:u _ | _ 178 _ | _ o:w:o _ | _ 199 _ | _ i:w:i _ | _ 102 _ | _ e:w:e _ | _ 190 _ | _ a:w:a _ | _ 149 _ | _ e:w:e _ | _ 169 _ | _ i:w:i _ | _ 186 _ | _ o:w:o _ | _ 00000000 _ | _ e.a.e.i. _ | _ 00000000 _ | _ 150 _ | _ u:w:u _ | _ 170 _ | _ o:w:o _ | _ 192 _ | _ i:w:i _ | _ 196 _ | _ e:w:e _ | _ 156 _ | _ a:w:a _ | _ 199 _ | _ e:w:e _ | _ 180 _ | _ i:w:i _ | _ 178 _ | _ o:w:o _ | _ 00000000 _ | _ u.o.i.e. _ | _ 00000000 _ | _ 151 _ | _ u:w:u _ | _ 170 _ | _ o:w:o _ | _ 191 _ | _ i:w:i _ | _ 196 _ | _ e:w:e _ | _ 182 _ | _ a:w:a _ | _ 141 _ | _ e:w:e _ | _ 161 _ | _ i:w:i _ | _ 178 _ | _ o:w:o _ | _ 00000000 _ | _ o.i.e.a. _ | _ 00000000 _ | _ 142 _ | _ u:w:u _ | _ 162 _ | _ o:w:o _ | _ 184 _ | _ i:w:i _ | _ 188 _ | _ e:w:e _ | _ 148 _ | _ a:w:a _ | _ 191 _ | _ e:w:e _ | _ 172 _ | _ i:w:i _ | _ 171 _ | _ o:w:o _ | _ 00000000 _ | _ i.e.a.e. _ | _ 00000000 _ | _ 143 _ | _ u:w:u _ | _ 162 _ | _ o:w:o _ | _ 183 _ | _ i:w:i _ | _ 188 _ | _ e:w:e _ | _ 174 _ | _ a:w:a _ | _ 133 _ | _ e:w:e _ | _ 153 _ | _ i:w:i _ | _ 171 _ | _ o:w:o _ | _ 00000000 _ | _ e.a.e.i. _ | _ 00000000 _ | _ 134 _ | _ u:w:u _ | _ 154 _ | _ o:w:o _ | _ 176 _ | _ i:w:i _ | _ 180 _ | _ e:w:e _ | _ 140 _ | _ a:w:a _ | _ 183 _ | _ e:w:e _ | _ 164 _ | _ i:w:i _ | _ 163 _ | _ o:w:o _ | _ 00000000 _ | _ u.o.i.e. _ | _ 00000000 _ | _ 135 _ | _ u:w:u _ | _ 154 _ | _ o:w:o _ | _ 175 _ | _ i:w:i _ | _ 180 _ | _ e:w:e _ | _ 166 _ | _ a:w:a _ | _ 125 _ | _ e:w:e _ | _ 145 _ | _ i:w:i _ | _ 163 _ | _ o:w:o _ | _ 00000000 _ | _ o.i.e.a. _ | _ 00000000 _ | _ 126 _ | _ u:w:u _ | _ 146 _ | _ o:w:o _ | _ 168 _ | _ i:w:i _ | _ 172 _ | _ e:w:e _ | _ 132 _ | _ a:w:a _ | _ 175 _ | _ e:w:e _ | _ 156 _ | _ i:w:i _ | _ 155 _ | _ o:w:o _ | _ 00000000 _ | _ i.e.a.e. _ | _ 00000000 _ | _ 127 _ | _ u:w:u _ | _ 146 _ | _ o:w:o _ | _ 167 _ | _ i:w:i _ | _ 172 _ | _ e:w:e _ | _ 158 _ | _ a:w:a _ | _ 117 _ | _ e:w:e _ | _ 137 _ | _ i:w:i _ | _ 155 _ | _ o:w:o _ | _ 00000000 _ | _ e.a.e.i. _ | _ 00000000 _ | _ 118 _ | _ u:w:u _ | _ 138 _ | _ o:w:o _ | _ 160 _ | _ i:w:i _ | _ 164 _ | _ e:w:e _ | _ 124 _ | _ a:w:a _ | _ 167 _ | _ e:w:e _ | _ 148 _ | _ i:w:i _ | _ 147 _ | _ o:w:o _ | _ 00000000 _ | _ u.o.i.e. _ | _ 00000000 _ | _ 119 _ | _ u:w:u _ | _ 138 _ | _ o:w:o _ | _ 159 _ | _ i:w:i _ | _ 164 _ | _ e:w:e _ | _ 150 _ | _ a:w:a _ | _ 109 _ | _ e:w:e _ | _ 129 _ | _ i:w:i _ | _ 147 _ | _ o:w:o _ | _ 00000000 _ | _ o.i.e.a. _ | _ 00000000 _ | _ 110 _ | _ u:w:u _ | _ 130 _ | _ o:w:o _ | _ 151 _ | _ i:w:i _ | _ 156 _ | _ e:w:e _ | _ 116 _ | _ a:w:a _ | _ 159 _ | _ e:w:e _ | _ 140 _ | _ i:w:i _ | _ 139 _ | _ o:w:o _ | _ 00000000 _ | _ i.e.a.e. _ | _ 00000000 _ | _ 111 _ | _ u:w:u _ | _ 130 _ | _ o:w:o _ | _ 151 _ | _ i:w:i _ | _ 156 _ | _ e:w:e _ | _ 142 _ | _ a:w:a _ | _ 101 _ | _ e:w:e _ | _ 121 _ | _ i:w:i _ | _ 139 _ | _ o:w:o _ | _ 00000000 _ | _ e.a.e.i. _ | _ 00000000 _ | _ 102 _ | _ u:w:u _ | _ 122 _ | _ o:w:o _ | _ 143 _ | _ i:w:i _ | _ 148 _ | _ e:w:e _ | _ 108 _ | _ a:w:a _ | _ 151 _ | _ e:w:e _ | _ 132 _ | _ i:w:i _ | _ 131 _ | _ o:w:o _ | _ 00000000 _ | _ u.o.i.e. _ | _ 00000000 _ | _ 103 _ | _ u:w:u _ | _ 122 _ | _ o:w:o _ | _ 143 _ | _ i:w:i _ | _ 148 _ | _ e:w:e _ | _ 134 _ | _ a:w:a _ | _ 193 _ | _ e:w:e _ | _ 113 _ | _ i:w:i _ | _ 131 _ | _ o:w:o _ | _ 00000000 _ | _ o.i.e.a. _ | _ 00000000 _ | _ 94 _ | _ u:w:u _ | _ 114 _ | _ o:w:o _ | _ 135 _ | _ i:w:i _ | _ 140 _ | _ e:w:e _ | _ 100 _ | _ a:w:a _ | _ 143 _ | _ e:w:e _ | _ 124 _ | _ i:w:i _ | _ 123 _ | _ o:w:o _ | _ 00000000 _ | _ i.e.a.e. _ | _ 00000000 _ | _ 95 _ | _ u:w:u _ | _ 114 _ | _ o:w:o _ | _ 135 _ | _ i:w:i _ | _ 140 _ | _ e:w:e _ | _ 126 _ | _ a:w:a _ | _ 185 _ | _ e:w:e _ | _ 105 _ | _ i:w:i _ | _ 123 _ | _ o:w:o _ | _ 00000000 _ | _ e.a.e.i. _ | _ 00000000 _ | _ 86 _ | _ u:w:u _ | _ 106 _ | _ o:w:o _ | _ 127 _ | _ i:w:i _ | _ 132 _ | _ e:w:e _ | _ 92 _ | _ a:w:a _ | _ 135 _ | _ e:w:e _ | _ 116 _ | _ i:w:i _ | _ 115 _ | _ o:w:o _ | _ 00000000 _ | _ u.o.i.e. _ | _ 00000000 _ | _ 83 _ | _ u:w:u _ | _ 106 _ | _ o:w:o _ | _ 127 _ | _ i:w:i _ | _ 132 _ | _ e:w:e _ | _ 118 _ | _ a:w:a _ | _ 177 _ | _ e:w:e _ | _ 97 _ | _ i:w:i _ | _ 115 _ | _ o:w:o _ | _ 00000000 _ | _ o.i.e.a. _ | _ 00000000 _ | _ 78 _ | _ u:w:u _ | _ 98 _ | _ o:w:o _ | _ 119 _ | _ i:w:i _ | _ 124 _ | _ e:w:e _ | _ 84 _ | _ a:w:a _ | _ 127 _ | _ e:w:e _ | _ 108 _ | _ i:w:i _ | _ 107 _ | _ o:w:o _ | _ 00000000 _ | _ i.e.a.e. _ | _ 00000000 _ | _ 75 _ | _ u:w:u _ | _ 98 _ | _ o:w:o _ | _ 119 _ | _ i:w:i _ | _ 124 _ | _ e:w:e _ | _ 110 _ | _ a:w:a _ | _ 169 _ | _ e:w:e _ | _ 89 _ | _ i:w:i _ | _ 107 _ | _ o:w:o _ | _ 00000000 _ | _ e.a.e.i. _ | _ 00000000 _ | _ 70 _ | _ u:w:u _ | _ 90 _ | _ o:w:o _ | _ 111 _ | _ i:w:i _ | _ 116 _ | _ e:w:e _ | _ 76 _ | _ a:w:a _ | _ 119 _ | _ e:w:e _ | _ 100 _ | _ i:w:i _ | _ 99 _ | _ o:w:o _ | _ 00000000 _ | _ u.o.i.e. _ | _ 00000000 _ | _ 67 _ | _ u:w:u _ | _ 90 _ | _ o:w:o _ | _ 111 _ | _ i:w:i _ | _ 116 _ | _ e:w:e _ | _ 102 _ | _ a:w:a _ | _ 161 _ | _ e:w:e _ | _ 81 _ | _ i:w:i _ | _ 99 _ | _ o:w:o _ | _ 00000000 _ | _ o.i.e.a. _ | _ 00000000 _ | _ 62 _ | _ u:w:u _ | _ 82 _ | _ o:w:o _ | _ 103 _ | _ i:w:i _ | _ 108 _ | _ e:w:e _ | _ 68 _ | _ a:w:a _ | _ 111 _ | _ e:w:e _ | _92_ | _ i:w:i _ | _ 91 _ | _ o:w:o _ | _ 00000000 _ | _ i.e.a.e. _ | _ 00000000 _ | _ 59 _ | _ u:w:u _ | _ 82 _ | _ o:w:o _ | _ 103 _ | _ i:w:i _ | _ 108 _ | _ e:w:e _ | _ 94 _ | _ a:w:a _ | _ 153 _ | _ e:w:e _ | _ 73 _ | _ i:w:i _ | _ 91 _ | _ o:w:o _ | _ 00000000 _ | _ e.a.e.i. _ | _ 00000000 _ | _ 54 _ | _ u:w:u _ | _ 74 _ | _ o:w:o _ | _ 95 _ | _ i:w:i _ | _ 100 _ | _ e:w:e _ | _ 60 _ | _ a:w:a _ | _ 103 _ | _ e:w:e _ | _ 84 _ | _ i:w:i _ | _ 83 _ | _ o:w:o _ | _ 00000000 _ | _ u.o.i.e. _ | _ 00000000 _ | _ 51 _ | _ u:w:u _ | _ 74 _ | _ o:w:o _ | _ 95 _ | _ i:w:i _ | _ 100 _ | _ e:w:e _ | _ 86 _ | _ a:w:a _ | _ 145 _ | _ e:w:e _ | _ 65 _ | _ i:w:i _ | _ 83 _ | _ o:w:o _ | _ 00000000 _ | _ o.i.e.a. _ | _ 00000000 _ | _ 46 _ | _ u:w:u _ | _ 66 _ | _ o:w:o _ | _ 87 _ | _ i:w:i _ | _ 92 _ | _ e:w:e _ | _ 52 _ | _ a:w:a _ | _ 95 _ | _ e:w:e _ | _ 76 _ | _ i:w:i _ | _ 75 _ | _ o:w:o _ | _ 00000000 _ | _ i.e.a.e. _ | _ 00000000 _ | _ 43_ | _ u:w:u _ | _ 66 _ | _ o:w:o _ | _ 87 _ | _ i:w:i _ | _ 92 _ | _ e:w:e _ | _ 78 _ | _ a:w:a _ | _ 137 _ | _ e:w:e _ | _ 57 _ | _ i:w:i _ | _ 75 _ | _ o:w:o _ | _ 00000000 _ | _ e.a.e.i. _ | _ 00000000 _ | _ 38 _ | _ u:w:u _ | _ 58 _ | _ o:w:o _ | _ 79 _ | _ i:w:i _ | _ 84 _ | _ e:w:e _ | _ 44 _ | _ a:w:a _ | _ 87 _ | _ e:w:e _ | _ 68 _ | _ i:w:i _ | _ 67 _ | _ o:w:o _ | _ 00000000 _ | _ u.o.i.e. _ | _ 00000000 _ | _ 35 _ | _ u:w:u _ | _ 58 _ | _ o:w:o _ | _ 79 _ | _ i:w:i _ | _ 84 _ | _ e:w:e _ | _ 70 _ | _ a:w:a _ | _ 129 _ | _ e:w:e _ | _ 49 _ | _ i:w:i _ | _ -67_ | _ o:w:o _ | _ 00000000 _ | _ o.i.e.a. _ | _ 00000000 _ | _ 30 _ | _ u:w:u _ | _ 50 _ | _ o:w:o _ | _ 71 _ | _ i:w:i _ | _ 76 _ | _ e:w:e _ | _ 36 _ | _ a:w:a _ | _ 79 _ | _ e:w:e _ | _ 60 _ | _ i:w:i _ | _ 59 _ | _ o:w:o _ | _ 00000000 _ | _ i.e.a.e. _ | _ 00000000 _ | _ 37 _ | _ u:w:u _ | _ 50 _ | _ o:w:o _ | _ 71 _ | _ i:w:i _ | _ 76 _ | _ e:w:e _ | _ 62 _ | _ a:w:a _ | _ 121 _ | _ e:w:e _ | _ 41 _ | _ i:w:i _ | _ 59 _ | _ o:w:o _ | _ 00000000 _ | _ e.a.e.i. _ | _ 00000000 _ | _ 22 _ | _ u:w:u _ | _ 42 _ | _ o:w:o _ | _ 63 _ | _ i:w:i _ | _ 68 _ | _ e:w:e _ | _ 28 _ | _ a:w:a _ | _ 71 _ | _ e:w:e _ | _ 52 _ | _ i:w:i _ | _ 51 _ | _ o:w:o _ | _ 00000000 _ | _ u.o.i.e. _ | _ 00000000 _ | _ 19 _ | _ u:w:u _ | _ 42 _ | _ o:w:o _ | _ 63 _ | _ i:w:i _ | _ 68 _ | _ e:w:e _ | _ 54 _ | _ a:w:a _ | _ 113 _ | _ e:w:e _ | _ 33 _ | _ i:w:i _ | _ 51 _ | _ o:w:o _ | _ 00000000 _ | _ o.i.e.a. _ | _ 00000000 _ | _ 14 _ | _ u:w:u _ | _ 34 _ | _ o:w:o _ | _ 55 _ | _ i:w:i _ | _ 60 _ | _ e:w:e _ | _ 20 _ | _ a:w:a _ | _ 63 _ | _ e:w:e _ | _ 44 _ | _ i:w:i _ | _ 43 _ | _ o:w:o _ | _ 00000000 _ | _ i.e.a.e. _ | _ 00000000 _ | _ 11 _ | _ u:w:u _ | _ 34 _ | _ o:w:o _ | _ 55 _ | _ i:w:i _ | _ 60 _ | _ e:w:e _ | _ 46 _ | _ a:w:a _ | _ 105 _ | _ e:w:e _ | _ 25 _ | _ i:w:i _ | _ 43 _ | _ o:w:o _ | _ 00000000 _ | _ e.a.e.i. _ | _ 00000000 _ | _ | _ 009-009-1963 _ ||